`timescale 1ns / 1ps


module tb_fourbitcla_claudehigh(

    );
endmodule
